package user_types is
    constant STREAM_SIZE : integer := 16;
end package user_types;